library ieee;
use ieee.std_logic_1164.all;

library work;

entity flipFlop_tb is
end;

architecture behaviour of flipFlop_tb is

signal clk_tb, clkEnable_tb, D_tb, Q_tb : std_logic;

component flipFlop is
   port(
      clk			: in std_logic;
      clkEnable	: in std_logic;
      D 				: in std_logic;
      Q				: out std_logic
   );
end component;

 
begin
	DUT1 : flipFlop port map(
		clk	=> clk_tb,
		clkEnable => clkEnable_tb,
		D => D_tb,
		Q => Q_tb	
	);
	
	sim_process: process
	begin
	
		wait for 1 ns;
		clk_tb		<= '0';
		clkEnable_tb		<= '1';
		D_tb<= '0';		
		wait for 9 ns;
		clk_tb		<= '1';
		wait for 10 ns;	
		clk_tb		<= '0';	
		wait for 10 ns;
		clk_tb		<= '1';
		D_tb <= '1';
		wait for 10 ns;		
		wait;
	end process sim_process;
end behaviour;