increment_inst : increment PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
