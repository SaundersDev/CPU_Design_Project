LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY regPC IS
	PORT(
		clk, clr, Rin : IN STD_LOGIC;
		BusMuxOut : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		BusMuxIn : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
END ENTITY regPC;

ARCHITECTURE arc OF regPC IS
BEGIN
	SingleRegister:
	PROCESS (clk, clr, Rin, BusMuxOut)
	BEGIN
		IF (clr = '0') THEN
			BusMuxIn <= (others => '0' );
		Elsif ((clr = '0') and rising_edge(clk) AND (Rin = '1')) THEN
			BusMuxIn <= BusMuxOut;
		END IF;
	END PROCESS;
END ARCHITECTURE arc;
